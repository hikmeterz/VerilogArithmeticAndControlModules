`timescale 1ns / 1ps
// Create Date: 13.11.2021 19:32:57


module bir_sayma(
    



    );
endmodule
